magic
tech scmos
timestamp 1732166173
<< error_p >>
rect 148 -561 149 -554
rect 175 -561 176 -554
rect 296 -601 297 -594
rect 291 -633 292 -630
rect 294 -637 295 -633
rect 148 -711 149 -704
rect 175 -711 176 -704
rect 296 -771 297 -764
rect 291 -803 292 -800
rect 294 -807 295 -803
rect 524 -851 525 -844
rect 624 -851 625 -844
rect 724 -851 725 -844
rect 824 -851 825 -844
rect 148 -861 149 -854
rect 175 -861 176 -854
rect 506 -895 507 -888
rect 606 -895 607 -888
rect 706 -895 707 -888
rect 806 -895 807 -888
rect 296 -941 297 -934
rect 291 -973 292 -970
rect 294 -977 295 -973
rect 148 -1011 149 -1004
rect 175 -1011 176 -1004
rect 296 -1111 297 -1104
rect 291 -1143 292 -1140
rect 294 -1147 295 -1143
<< nwell >>
rect 228 -525 339 -496
rect 5 -589 120 -526
rect 300 -549 325 -525
rect 5 -739 120 -676
rect 228 -695 339 -666
rect 300 -719 325 -695
rect 5 -889 120 -826
rect 463 -834 502 -813
rect 228 -865 339 -836
rect 511 -845 534 -818
rect 563 -834 602 -813
rect 611 -845 634 -818
rect 663 -834 702 -813
rect 711 -845 734 -818
rect 763 -834 802 -813
rect 811 -845 834 -818
rect 300 -889 325 -865
rect 5 -1039 120 -976
rect 228 -1035 339 -1006
rect 300 -1059 325 -1035
<< polysilicon >>
rect 238 -513 246 -511
rect 266 -513 272 -511
rect 294 -513 300 -511
rect 320 -513 328 -511
rect 311 -523 313 -520
rect 145 -533 147 -530
rect 172 -533 174 -530
rect 15 -545 25 -543
rect 45 -545 54 -543
rect 69 -545 82 -543
rect 102 -545 109 -543
rect 145 -557 147 -553
rect 172 -557 174 -553
rect 146 -561 147 -557
rect 173 -561 174 -557
rect 311 -560 313 -543
rect 145 -565 147 -561
rect 172 -565 174 -561
rect 15 -570 25 -568
rect 45 -570 52 -568
rect 72 -570 82 -568
rect 102 -570 109 -568
rect 311 -574 313 -570
rect 145 -579 147 -575
rect 172 -579 174 -575
rect 293 -584 295 -580
rect 293 -597 295 -594
rect 13 -603 29 -601
rect 39 -603 47 -601
rect 74 -603 86 -601
rect 96 -603 105 -601
rect 294 -600 295 -597
rect 293 -617 295 -613
rect 14 -633 29 -631
rect 39 -633 50 -631
rect 77 -633 86 -631
rect 96 -633 105 -631
rect 293 -633 295 -627
rect 293 -637 294 -633
rect 145 -683 147 -680
rect 172 -683 174 -680
rect 15 -695 25 -693
rect 45 -695 54 -693
rect 69 -695 82 -693
rect 102 -695 109 -693
rect 238 -683 246 -681
rect 266 -683 272 -681
rect 294 -683 300 -681
rect 320 -683 328 -681
rect 311 -693 313 -690
rect 145 -707 147 -703
rect 172 -707 174 -703
rect 146 -711 147 -707
rect 173 -711 174 -707
rect 145 -715 147 -711
rect 172 -715 174 -711
rect 15 -720 25 -718
rect 45 -720 52 -718
rect 72 -720 82 -718
rect 102 -720 109 -718
rect 145 -729 147 -725
rect 172 -729 174 -725
rect 311 -730 313 -713
rect 311 -744 313 -740
rect 13 -753 29 -751
rect 39 -753 47 -751
rect 74 -753 86 -751
rect 96 -753 105 -751
rect 293 -754 295 -750
rect 293 -767 295 -764
rect 294 -770 295 -767
rect 14 -783 29 -781
rect 39 -783 50 -781
rect 77 -783 86 -781
rect 96 -783 105 -781
rect 293 -787 295 -783
rect 293 -803 295 -797
rect 293 -807 294 -803
rect 521 -823 523 -821
rect 621 -823 623 -821
rect 721 -823 723 -821
rect 821 -823 823 -821
rect 473 -826 476 -824
rect 496 -826 505 -824
rect 145 -833 147 -830
rect 172 -833 174 -830
rect 15 -845 25 -843
rect 45 -845 54 -843
rect 69 -845 82 -843
rect 102 -845 109 -843
rect 483 -842 485 -839
rect 145 -857 147 -853
rect 172 -857 174 -853
rect 238 -853 246 -851
rect 266 -853 272 -851
rect 294 -853 300 -851
rect 320 -853 328 -851
rect 146 -861 147 -857
rect 173 -861 174 -857
rect 573 -826 576 -824
rect 596 -826 605 -824
rect 583 -842 585 -839
rect 521 -847 523 -843
rect 522 -851 523 -847
rect 483 -855 485 -852
rect 521 -854 523 -851
rect 673 -826 676 -824
rect 696 -826 705 -824
rect 683 -842 685 -839
rect 621 -847 623 -843
rect 622 -851 623 -847
rect 503 -858 505 -855
rect 145 -865 147 -861
rect 172 -865 174 -861
rect 311 -863 313 -860
rect 15 -870 25 -868
rect 45 -870 52 -868
rect 72 -870 82 -868
rect 102 -870 109 -868
rect 145 -879 147 -875
rect 172 -879 174 -875
rect 583 -855 585 -852
rect 621 -854 623 -851
rect 773 -826 776 -824
rect 796 -826 805 -824
rect 783 -842 785 -839
rect 721 -847 723 -843
rect 722 -851 723 -847
rect 603 -858 605 -855
rect 503 -877 505 -868
rect 521 -869 523 -864
rect 683 -855 685 -852
rect 721 -854 723 -851
rect 821 -847 823 -843
rect 822 -851 823 -847
rect 703 -858 705 -855
rect 603 -877 605 -868
rect 621 -869 623 -864
rect 783 -855 785 -852
rect 821 -854 823 -851
rect 803 -858 805 -855
rect 703 -877 705 -868
rect 721 -869 723 -864
rect 803 -877 805 -868
rect 821 -869 823 -864
rect 311 -900 313 -883
rect 504 -895 505 -891
rect 604 -895 605 -891
rect 704 -895 705 -891
rect 804 -895 805 -891
rect 503 -899 505 -895
rect 603 -899 605 -895
rect 703 -899 705 -895
rect 803 -899 805 -895
rect 13 -903 29 -901
rect 39 -903 47 -901
rect 74 -903 86 -901
rect 96 -903 105 -901
rect 311 -914 313 -910
rect 503 -912 505 -909
rect 603 -912 605 -909
rect 703 -912 705 -909
rect 803 -912 805 -909
rect 293 -924 295 -920
rect 14 -933 29 -931
rect 39 -933 50 -931
rect 77 -933 86 -931
rect 96 -933 105 -931
rect 293 -937 295 -934
rect 294 -940 295 -937
rect 293 -957 295 -953
rect 293 -973 295 -967
rect 293 -977 294 -973
rect 145 -983 147 -980
rect 172 -983 174 -980
rect 15 -995 25 -993
rect 45 -995 54 -993
rect 69 -995 82 -993
rect 102 -995 109 -993
rect 145 -1007 147 -1003
rect 172 -1007 174 -1003
rect 146 -1011 147 -1007
rect 173 -1011 174 -1007
rect 145 -1015 147 -1011
rect 172 -1015 174 -1011
rect 15 -1020 25 -1018
rect 45 -1020 52 -1018
rect 72 -1020 82 -1018
rect 102 -1020 109 -1018
rect 238 -1023 246 -1021
rect 266 -1023 272 -1021
rect 294 -1023 300 -1021
rect 320 -1023 328 -1021
rect 145 -1029 147 -1025
rect 172 -1029 174 -1025
rect 311 -1033 313 -1030
rect 13 -1053 29 -1051
rect 39 -1053 47 -1051
rect 74 -1053 86 -1051
rect 96 -1053 105 -1051
rect 311 -1070 313 -1053
rect 14 -1083 29 -1081
rect 39 -1083 50 -1081
rect 77 -1083 86 -1081
rect 96 -1083 105 -1081
rect 311 -1084 313 -1080
rect 293 -1094 295 -1090
rect 293 -1107 295 -1104
rect 294 -1110 295 -1107
rect 293 -1127 295 -1123
rect 293 -1143 295 -1137
rect 293 -1147 294 -1143
<< ndiffusion >>
rect 144 -575 145 -565
rect 147 -575 148 -565
rect 171 -575 172 -565
rect 174 -575 175 -565
rect 310 -570 311 -560
rect 313 -570 314 -560
rect 292 -594 293 -584
rect 295 -594 296 -584
rect 29 -601 39 -600
rect 86 -601 96 -600
rect 29 -604 39 -603
rect 86 -604 96 -603
rect 29 -631 39 -630
rect 292 -627 293 -617
rect 295 -627 296 -617
rect 86 -631 96 -630
rect 29 -634 39 -633
rect 86 -634 96 -633
rect 144 -725 145 -715
rect 147 -725 148 -715
rect 171 -725 172 -715
rect 174 -725 175 -715
rect 310 -740 311 -730
rect 313 -740 314 -730
rect 29 -751 39 -750
rect 86 -751 96 -750
rect 29 -754 39 -753
rect 86 -754 96 -753
rect 292 -764 293 -754
rect 295 -764 296 -754
rect 29 -781 39 -780
rect 86 -781 96 -780
rect 29 -784 39 -783
rect 86 -784 96 -783
rect 292 -797 293 -787
rect 295 -797 296 -787
rect 482 -852 483 -842
rect 485 -852 486 -842
rect 582 -852 583 -842
rect 585 -852 586 -842
rect 144 -875 145 -865
rect 147 -875 148 -865
rect 171 -875 172 -865
rect 174 -875 175 -865
rect 502 -868 503 -858
rect 505 -868 506 -858
rect 520 -864 521 -854
rect 523 -864 524 -854
rect 682 -852 683 -842
rect 685 -852 686 -842
rect 602 -868 603 -858
rect 605 -868 606 -858
rect 620 -864 621 -854
rect 623 -864 624 -854
rect 782 -852 783 -842
rect 785 -852 786 -842
rect 702 -868 703 -858
rect 705 -868 706 -858
rect 720 -864 721 -854
rect 723 -864 724 -854
rect 802 -868 803 -858
rect 805 -868 806 -858
rect 820 -864 821 -854
rect 823 -864 824 -854
rect 29 -901 39 -900
rect 86 -901 96 -900
rect 29 -904 39 -903
rect 86 -904 96 -903
rect 310 -910 311 -900
rect 313 -910 314 -900
rect 502 -909 503 -899
rect 505 -909 506 -899
rect 602 -909 603 -899
rect 605 -909 606 -899
rect 702 -909 703 -899
rect 705 -909 706 -899
rect 802 -909 803 -899
rect 805 -909 806 -899
rect 29 -931 39 -930
rect 86 -931 96 -930
rect 29 -934 39 -933
rect 86 -934 96 -933
rect 292 -934 293 -924
rect 295 -934 296 -924
rect 292 -967 293 -957
rect 295 -967 296 -957
rect 144 -1025 145 -1015
rect 147 -1025 148 -1015
rect 171 -1025 172 -1015
rect 174 -1025 175 -1015
rect 29 -1051 39 -1050
rect 86 -1051 96 -1050
rect 29 -1054 39 -1053
rect 86 -1054 96 -1053
rect 29 -1081 39 -1080
rect 310 -1080 311 -1070
rect 313 -1080 314 -1070
rect 86 -1081 96 -1080
rect 29 -1084 39 -1083
rect 86 -1084 96 -1083
rect 292 -1104 293 -1094
rect 295 -1104 296 -1094
rect 292 -1137 293 -1127
rect 295 -1137 296 -1127
<< pdiffusion >>
rect 246 -511 266 -510
rect 300 -511 320 -510
rect 246 -514 266 -513
rect 300 -514 320 -513
rect 25 -543 45 -542
rect 82 -543 102 -542
rect 25 -546 45 -545
rect 82 -546 102 -545
rect 144 -553 145 -533
rect 147 -553 148 -533
rect 171 -553 172 -533
rect 174 -553 175 -533
rect 310 -543 311 -523
rect 313 -543 314 -523
rect 25 -568 45 -567
rect 82 -568 102 -567
rect 25 -571 45 -570
rect 82 -571 102 -570
rect 25 -693 45 -692
rect 82 -693 102 -692
rect 25 -696 45 -695
rect 82 -696 102 -695
rect 144 -703 145 -683
rect 147 -703 148 -683
rect 171 -703 172 -683
rect 174 -703 175 -683
rect 246 -681 266 -680
rect 300 -681 320 -680
rect 246 -684 266 -683
rect 300 -684 320 -683
rect 25 -718 45 -717
rect 310 -713 311 -693
rect 313 -713 314 -693
rect 82 -718 102 -717
rect 25 -721 45 -720
rect 82 -721 102 -720
rect 476 -824 496 -823
rect 476 -827 496 -826
rect 25 -843 45 -842
rect 82 -843 102 -842
rect 25 -846 45 -845
rect 82 -846 102 -845
rect 144 -853 145 -833
rect 147 -853 148 -833
rect 171 -853 172 -833
rect 174 -853 175 -833
rect 246 -851 266 -850
rect 300 -851 320 -850
rect 246 -854 266 -853
rect 300 -854 320 -853
rect 520 -843 521 -823
rect 523 -843 524 -823
rect 576 -824 596 -823
rect 576 -827 596 -826
rect 620 -843 621 -823
rect 623 -843 624 -823
rect 676 -824 696 -823
rect 676 -827 696 -826
rect 25 -868 45 -867
rect 82 -868 102 -867
rect 25 -871 45 -870
rect 82 -871 102 -870
rect 310 -883 311 -863
rect 313 -883 314 -863
rect 720 -843 721 -823
rect 723 -843 724 -823
rect 776 -824 796 -823
rect 776 -827 796 -826
rect 820 -843 821 -823
rect 823 -843 824 -823
rect 25 -993 45 -992
rect 82 -993 102 -992
rect 25 -996 45 -995
rect 82 -996 102 -995
rect 144 -1003 145 -983
rect 147 -1003 148 -983
rect 171 -1003 172 -983
rect 174 -1003 175 -983
rect 25 -1018 45 -1017
rect 82 -1018 102 -1017
rect 25 -1021 45 -1020
rect 82 -1021 102 -1020
rect 246 -1021 266 -1020
rect 300 -1021 320 -1020
rect 246 -1024 266 -1023
rect 300 -1024 320 -1023
rect 310 -1053 311 -1033
rect 313 -1053 314 -1033
<< metal1 >>
rect 266 -510 300 -506
rect 332 -514 333 -510
rect 21 -528 82 -524
rect 21 -542 25 -528
rect 78 -542 82 -528
rect 138 -529 150 -525
rect 165 -529 177 -525
rect 140 -533 144 -529
rect 167 -533 171 -529
rect 2 -546 11 -542
rect 113 -546 122 -542
rect 45 -567 49 -546
rect 102 -567 106 -546
rect 136 -561 142 -557
rect 148 -565 152 -553
rect 164 -561 169 -557
rect 175 -565 179 -553
rect 2 -571 11 -567
rect 113 -571 122 -567
rect 21 -585 25 -571
rect 78 -585 82 -571
rect 140 -582 144 -575
rect 167 -582 171 -575
rect 137 -585 148 -582
rect 164 -585 175 -582
rect 21 -589 89 -585
rect 21 -596 25 -589
rect 78 -596 82 -589
rect 21 -600 29 -596
rect 78 -600 86 -596
rect 234 -597 238 -514
rect 266 -518 300 -514
rect 288 -552 292 -518
rect 306 -547 310 -543
rect 288 -556 306 -552
rect 288 -584 292 -556
rect 314 -560 318 -543
rect 306 -574 310 -570
rect 300 -594 301 -584
rect 0 -604 9 -600
rect 109 -604 118 -600
rect 234 -601 289 -597
rect 39 -630 43 -604
rect 96 -630 100 -604
rect 296 -617 301 -594
rect 300 -627 301 -617
rect 1 -634 10 -630
rect 109 -634 118 -630
rect 39 -645 43 -634
rect 96 -645 100 -634
rect 288 -643 292 -627
rect 328 -633 333 -514
rect 298 -637 333 -633
rect 39 -649 100 -645
rect 276 -647 305 -643
rect 21 -678 82 -674
rect 21 -692 25 -678
rect 78 -692 82 -678
rect 138 -679 150 -675
rect 165 -679 177 -675
rect 140 -683 144 -679
rect 167 -683 171 -679
rect 266 -680 300 -676
rect 2 -696 11 -692
rect 113 -696 122 -692
rect 45 -717 49 -696
rect 102 -717 106 -696
rect 136 -711 142 -707
rect 148 -715 152 -703
rect 164 -711 169 -707
rect 175 -715 179 -703
rect 2 -721 11 -717
rect 113 -721 122 -717
rect 21 -735 25 -721
rect 78 -735 82 -721
rect 332 -684 333 -680
rect 140 -732 144 -725
rect 167 -732 171 -725
rect 137 -735 148 -732
rect 164 -735 175 -732
rect 21 -739 89 -735
rect 21 -746 25 -739
rect 78 -746 82 -739
rect 21 -750 29 -746
rect 78 -750 86 -746
rect 0 -754 9 -750
rect 109 -754 118 -750
rect 39 -780 43 -754
rect 96 -780 100 -754
rect 234 -767 238 -684
rect 266 -688 300 -684
rect 288 -722 292 -688
rect 306 -717 310 -713
rect 288 -726 306 -722
rect 288 -754 292 -726
rect 314 -730 318 -713
rect 306 -744 310 -740
rect 300 -764 301 -754
rect 234 -771 289 -767
rect 1 -784 10 -780
rect 109 -784 118 -780
rect 39 -795 43 -784
rect 96 -795 100 -784
rect 296 -787 301 -764
rect 39 -799 100 -795
rect 300 -797 301 -787
rect 288 -813 292 -797
rect 328 -803 333 -684
rect 298 -807 333 -803
rect 276 -817 305 -813
rect 496 -823 520 -819
rect 596 -823 620 -819
rect 696 -823 720 -819
rect 796 -823 820 -819
rect 21 -828 82 -824
rect 21 -842 25 -828
rect 78 -842 82 -828
rect 138 -829 150 -825
rect 165 -829 177 -825
rect 464 -827 469 -823
rect 140 -833 144 -829
rect 167 -833 171 -829
rect 496 -831 502 -827
rect 2 -846 11 -842
rect 113 -846 122 -842
rect 45 -867 49 -846
rect 102 -867 106 -846
rect 479 -839 482 -835
rect 266 -850 300 -846
rect 136 -861 142 -857
rect 148 -865 152 -853
rect 164 -861 169 -857
rect 175 -865 179 -853
rect 2 -871 11 -867
rect 113 -871 122 -867
rect 21 -885 25 -871
rect 78 -885 82 -871
rect 332 -854 333 -850
rect 140 -882 144 -875
rect 167 -882 171 -875
rect 137 -885 148 -882
rect 164 -885 175 -882
rect 21 -889 89 -885
rect 21 -896 25 -889
rect 78 -896 82 -889
rect 21 -900 29 -896
rect 78 -900 86 -896
rect 0 -904 9 -900
rect 109 -904 118 -900
rect 39 -930 43 -904
rect 96 -930 100 -904
rect 1 -934 10 -930
rect 109 -934 118 -930
rect 39 -945 43 -934
rect 96 -945 100 -934
rect 234 -937 238 -854
rect 266 -858 300 -854
rect 288 -892 292 -858
rect 306 -887 310 -883
rect 288 -896 306 -892
rect 288 -924 292 -896
rect 314 -900 318 -883
rect 306 -914 310 -910
rect 300 -934 301 -924
rect 234 -941 289 -937
rect 39 -949 100 -945
rect 296 -957 301 -934
rect 300 -967 301 -957
rect 21 -978 82 -974
rect 21 -992 25 -978
rect 78 -992 82 -978
rect 138 -979 150 -975
rect 165 -979 177 -975
rect 140 -983 144 -979
rect 167 -983 171 -979
rect 288 -983 292 -967
rect 328 -973 333 -854
rect 478 -856 482 -852
rect 498 -847 502 -831
rect 564 -827 569 -823
rect 596 -831 602 -827
rect 579 -839 582 -835
rect 498 -851 518 -847
rect 498 -852 502 -851
rect 486 -856 502 -852
rect 524 -854 528 -843
rect 498 -858 502 -856
rect 492 -877 499 -873
rect 496 -895 500 -891
rect 506 -899 510 -868
rect 578 -856 582 -852
rect 598 -847 602 -831
rect 664 -827 669 -823
rect 696 -831 702 -827
rect 679 -839 682 -835
rect 598 -851 618 -847
rect 598 -852 602 -851
rect 586 -856 602 -852
rect 624 -854 628 -843
rect 598 -858 602 -856
rect 516 -869 520 -864
rect 592 -877 599 -873
rect 596 -895 600 -891
rect 606 -899 610 -868
rect 678 -856 682 -852
rect 698 -847 702 -831
rect 764 -827 769 -823
rect 796 -831 802 -827
rect 779 -839 782 -835
rect 698 -851 718 -847
rect 698 -852 702 -851
rect 686 -856 702 -852
rect 724 -854 728 -843
rect 698 -858 702 -856
rect 616 -869 620 -864
rect 692 -877 699 -873
rect 696 -895 700 -891
rect 706 -899 710 -868
rect 778 -856 782 -852
rect 798 -847 802 -831
rect 798 -851 818 -847
rect 798 -852 802 -851
rect 786 -856 802 -852
rect 824 -854 828 -843
rect 798 -858 802 -856
rect 716 -869 720 -864
rect 792 -877 799 -873
rect 796 -895 800 -891
rect 806 -899 810 -868
rect 816 -869 820 -864
rect 498 -913 502 -909
rect 598 -913 602 -909
rect 698 -913 702 -909
rect 798 -913 802 -909
rect 298 -977 333 -973
rect 2 -996 11 -992
rect 113 -996 122 -992
rect 45 -1017 49 -996
rect 102 -1017 106 -996
rect 276 -987 305 -983
rect 136 -1011 142 -1007
rect 148 -1015 152 -1003
rect 164 -1011 169 -1007
rect 175 -1015 179 -1003
rect 2 -1021 11 -1017
rect 113 -1021 122 -1017
rect 21 -1035 25 -1021
rect 78 -1035 82 -1021
rect 266 -1020 300 -1016
rect 332 -1024 333 -1020
rect 140 -1032 144 -1025
rect 167 -1032 171 -1025
rect 137 -1035 148 -1032
rect 164 -1035 175 -1032
rect 21 -1039 89 -1035
rect 21 -1046 25 -1039
rect 78 -1046 82 -1039
rect 21 -1050 29 -1046
rect 78 -1050 86 -1046
rect 0 -1054 9 -1050
rect 109 -1054 118 -1050
rect 39 -1080 43 -1054
rect 96 -1080 100 -1054
rect 1 -1084 10 -1080
rect 109 -1084 118 -1080
rect 39 -1095 43 -1084
rect 96 -1095 100 -1084
rect 39 -1099 100 -1095
rect 234 -1107 238 -1024
rect 266 -1028 300 -1024
rect 288 -1062 292 -1028
rect 306 -1057 310 -1053
rect 288 -1066 306 -1062
rect 288 -1094 292 -1066
rect 314 -1070 318 -1053
rect 306 -1084 310 -1080
rect 300 -1104 301 -1094
rect 234 -1111 289 -1107
rect 296 -1127 301 -1104
rect 300 -1137 301 -1127
rect 288 -1153 292 -1137
rect 328 -1143 333 -1024
rect 298 -1147 333 -1143
rect 276 -1157 305 -1153
<< ntransistor >>
rect 145 -575 147 -565
rect 172 -575 174 -565
rect 311 -570 313 -560
rect 293 -594 295 -584
rect 29 -603 39 -601
rect 86 -603 96 -601
rect 293 -627 295 -617
rect 29 -633 39 -631
rect 86 -633 96 -631
rect 145 -725 147 -715
rect 172 -725 174 -715
rect 311 -740 313 -730
rect 29 -753 39 -751
rect 86 -753 96 -751
rect 293 -764 295 -754
rect 29 -783 39 -781
rect 86 -783 96 -781
rect 293 -797 295 -787
rect 483 -852 485 -842
rect 583 -852 585 -842
rect 145 -875 147 -865
rect 172 -875 174 -865
rect 503 -868 505 -858
rect 521 -864 523 -854
rect 683 -852 685 -842
rect 603 -868 605 -858
rect 621 -864 623 -854
rect 783 -852 785 -842
rect 703 -868 705 -858
rect 721 -864 723 -854
rect 803 -868 805 -858
rect 821 -864 823 -854
rect 29 -903 39 -901
rect 86 -903 96 -901
rect 311 -910 313 -900
rect 503 -909 505 -899
rect 603 -909 605 -899
rect 703 -909 705 -899
rect 803 -909 805 -899
rect 29 -933 39 -931
rect 86 -933 96 -931
rect 293 -934 295 -924
rect 293 -967 295 -957
rect 145 -1025 147 -1015
rect 172 -1025 174 -1015
rect 29 -1053 39 -1051
rect 86 -1053 96 -1051
rect 311 -1080 313 -1070
rect 29 -1083 39 -1081
rect 86 -1083 96 -1081
rect 293 -1104 295 -1094
rect 293 -1137 295 -1127
<< ptransistor >>
rect 246 -513 266 -511
rect 300 -513 320 -511
rect 25 -545 45 -543
rect 82 -545 102 -543
rect 145 -553 147 -533
rect 172 -553 174 -533
rect 311 -543 313 -523
rect 25 -570 45 -568
rect 82 -570 102 -568
rect 25 -695 45 -693
rect 82 -695 102 -693
rect 145 -703 147 -683
rect 172 -703 174 -683
rect 246 -683 266 -681
rect 300 -683 320 -681
rect 311 -713 313 -693
rect 25 -720 45 -718
rect 82 -720 102 -718
rect 476 -826 496 -824
rect 25 -845 45 -843
rect 82 -845 102 -843
rect 145 -853 147 -833
rect 172 -853 174 -833
rect 246 -853 266 -851
rect 300 -853 320 -851
rect 521 -843 523 -823
rect 576 -826 596 -824
rect 621 -843 623 -823
rect 676 -826 696 -824
rect 25 -870 45 -868
rect 82 -870 102 -868
rect 311 -883 313 -863
rect 721 -843 723 -823
rect 776 -826 796 -824
rect 821 -843 823 -823
rect 25 -995 45 -993
rect 82 -995 102 -993
rect 145 -1003 147 -983
rect 172 -1003 174 -983
rect 25 -1020 45 -1018
rect 82 -1020 102 -1018
rect 246 -1023 266 -1021
rect 300 -1023 320 -1021
rect 311 -1053 313 -1033
<< polycontact >>
rect 234 -514 238 -510
rect 328 -514 332 -510
rect 11 -546 15 -542
rect 109 -546 113 -542
rect 306 -556 311 -552
rect 142 -561 146 -557
rect 169 -561 173 -557
rect 11 -571 15 -567
rect 109 -571 113 -567
rect 9 -604 13 -600
rect 105 -604 109 -600
rect 289 -601 294 -597
rect 10 -634 14 -630
rect 105 -634 109 -630
rect 294 -637 298 -633
rect 11 -696 15 -692
rect 109 -696 113 -692
rect 234 -684 238 -680
rect 328 -684 332 -680
rect 142 -711 146 -707
rect 169 -711 173 -707
rect 11 -721 15 -717
rect 109 -721 113 -717
rect 306 -726 311 -722
rect 9 -754 13 -750
rect 105 -754 109 -750
rect 289 -771 294 -767
rect 10 -784 14 -780
rect 105 -784 109 -780
rect 294 -807 298 -803
rect 469 -827 473 -823
rect 11 -846 15 -842
rect 109 -846 113 -842
rect 482 -839 486 -835
rect 234 -854 238 -850
rect 142 -861 146 -857
rect 169 -861 173 -857
rect 328 -854 332 -850
rect 569 -827 573 -823
rect 582 -839 586 -835
rect 518 -851 522 -847
rect 669 -827 673 -823
rect 682 -839 686 -835
rect 618 -851 622 -847
rect 11 -871 15 -867
rect 109 -871 113 -867
rect 769 -827 773 -823
rect 782 -839 786 -835
rect 718 -851 722 -847
rect 499 -877 503 -873
rect 818 -851 822 -847
rect 599 -877 603 -873
rect 699 -877 703 -873
rect 799 -877 803 -873
rect 306 -896 311 -892
rect 9 -904 13 -900
rect 500 -895 504 -891
rect 600 -895 604 -891
rect 700 -895 704 -891
rect 800 -895 804 -891
rect 105 -904 109 -900
rect 10 -934 14 -930
rect 105 -934 109 -930
rect 289 -941 294 -937
rect 294 -977 298 -973
rect 11 -996 15 -992
rect 109 -996 113 -992
rect 142 -1011 146 -1007
rect 169 -1011 173 -1007
rect 11 -1021 15 -1017
rect 109 -1021 113 -1017
rect 234 -1024 238 -1020
rect 328 -1024 332 -1020
rect 9 -1054 13 -1050
rect 105 -1054 109 -1050
rect 306 -1066 311 -1062
rect 10 -1084 14 -1080
rect 105 -1084 109 -1080
rect 289 -1111 294 -1107
rect 294 -1147 298 -1143
<< ndcontact >>
rect 140 -575 144 -565
rect 148 -575 152 -565
rect 167 -575 171 -565
rect 175 -575 179 -565
rect 306 -570 310 -560
rect 314 -570 318 -560
rect 288 -594 292 -584
rect 296 -594 300 -584
rect 29 -600 39 -596
rect 86 -600 96 -596
rect 29 -608 39 -604
rect 86 -608 96 -604
rect 29 -630 39 -626
rect 86 -630 96 -626
rect 288 -627 292 -617
rect 296 -627 300 -617
rect 29 -638 39 -634
rect 86 -638 96 -634
rect 140 -725 144 -715
rect 148 -725 152 -715
rect 167 -725 171 -715
rect 175 -725 179 -715
rect 306 -740 310 -730
rect 314 -740 318 -730
rect 29 -750 39 -746
rect 86 -750 96 -746
rect 29 -758 39 -754
rect 86 -758 96 -754
rect 288 -764 292 -754
rect 296 -764 300 -754
rect 29 -780 39 -776
rect 86 -780 96 -776
rect 29 -788 39 -784
rect 86 -788 96 -784
rect 288 -797 292 -787
rect 296 -797 300 -787
rect 478 -852 482 -842
rect 486 -852 490 -842
rect 578 -852 582 -842
rect 586 -852 590 -842
rect 140 -875 144 -865
rect 148 -875 152 -865
rect 167 -875 171 -865
rect 175 -875 179 -865
rect 498 -868 502 -858
rect 506 -868 510 -858
rect 516 -864 520 -854
rect 524 -864 528 -854
rect 678 -852 682 -842
rect 686 -852 690 -842
rect 598 -868 602 -858
rect 606 -868 610 -858
rect 616 -864 620 -854
rect 624 -864 628 -854
rect 778 -852 782 -842
rect 786 -852 790 -842
rect 698 -868 702 -858
rect 706 -868 710 -858
rect 716 -864 720 -854
rect 724 -864 728 -854
rect 798 -868 802 -858
rect 806 -868 810 -858
rect 816 -864 820 -854
rect 824 -864 828 -854
rect 29 -900 39 -896
rect 86 -900 96 -896
rect 29 -908 39 -904
rect 86 -908 96 -904
rect 306 -910 310 -900
rect 314 -910 318 -900
rect 498 -909 502 -899
rect 506 -909 510 -899
rect 598 -909 602 -899
rect 606 -909 610 -899
rect 698 -909 702 -899
rect 706 -909 710 -899
rect 798 -909 802 -899
rect 806 -909 810 -899
rect 29 -930 39 -926
rect 86 -930 96 -926
rect 29 -938 39 -934
rect 288 -934 292 -924
rect 296 -934 300 -924
rect 86 -938 96 -934
rect 288 -967 292 -957
rect 296 -967 300 -957
rect 140 -1025 144 -1015
rect 148 -1025 152 -1015
rect 167 -1025 171 -1015
rect 175 -1025 179 -1015
rect 29 -1050 39 -1046
rect 86 -1050 96 -1046
rect 29 -1058 39 -1054
rect 86 -1058 96 -1054
rect 29 -1080 39 -1076
rect 86 -1080 96 -1076
rect 306 -1080 310 -1070
rect 314 -1080 318 -1070
rect 29 -1088 39 -1084
rect 86 -1088 96 -1084
rect 288 -1104 292 -1094
rect 296 -1104 300 -1094
rect 288 -1137 292 -1127
rect 296 -1137 300 -1127
<< pdcontact >>
rect 246 -510 266 -506
rect 300 -510 320 -506
rect 246 -518 266 -514
rect 300 -518 320 -514
rect 25 -542 45 -538
rect 82 -542 102 -538
rect 25 -550 45 -546
rect 82 -550 102 -546
rect 140 -553 144 -533
rect 148 -553 152 -533
rect 167 -553 171 -533
rect 175 -553 179 -533
rect 306 -543 310 -523
rect 314 -543 318 -523
rect 25 -567 45 -563
rect 82 -567 102 -563
rect 25 -575 45 -571
rect 82 -575 102 -571
rect 246 -680 266 -676
rect 25 -692 45 -688
rect 82 -692 102 -688
rect 25 -700 45 -696
rect 82 -700 102 -696
rect 140 -703 144 -683
rect 148 -703 152 -683
rect 167 -703 171 -683
rect 175 -703 179 -683
rect 300 -680 320 -676
rect 246 -688 266 -684
rect 300 -688 320 -684
rect 25 -717 45 -713
rect 82 -717 102 -713
rect 306 -713 310 -693
rect 314 -713 318 -693
rect 25 -725 45 -721
rect 82 -725 102 -721
rect 476 -823 496 -819
rect 576 -823 596 -819
rect 676 -823 696 -819
rect 776 -823 796 -819
rect 476 -831 496 -827
rect 25 -842 45 -838
rect 82 -842 102 -838
rect 25 -850 45 -846
rect 82 -850 102 -846
rect 140 -853 144 -833
rect 148 -853 152 -833
rect 167 -853 171 -833
rect 175 -853 179 -833
rect 246 -850 266 -846
rect 300 -850 320 -846
rect 246 -858 266 -854
rect 516 -843 520 -823
rect 524 -843 528 -823
rect 576 -831 596 -827
rect 300 -858 320 -854
rect 616 -843 620 -823
rect 624 -843 628 -823
rect 676 -831 696 -827
rect 25 -867 45 -863
rect 82 -867 102 -863
rect 25 -875 45 -871
rect 82 -875 102 -871
rect 306 -883 310 -863
rect 314 -883 318 -863
rect 716 -843 720 -823
rect 724 -843 728 -823
rect 776 -831 796 -827
rect 816 -843 820 -823
rect 824 -843 828 -823
rect 25 -992 45 -988
rect 82 -992 102 -988
rect 25 -1000 45 -996
rect 82 -1000 102 -996
rect 140 -1003 144 -983
rect 148 -1003 152 -983
rect 167 -1003 171 -983
rect 175 -1003 179 -983
rect 25 -1017 45 -1013
rect 82 -1017 102 -1013
rect 25 -1025 45 -1021
rect 82 -1025 102 -1021
rect 246 -1020 266 -1016
rect 300 -1020 320 -1016
rect 246 -1028 266 -1024
rect 300 -1028 320 -1024
rect 306 -1053 310 -1033
rect 314 -1053 318 -1033
<< labels >>
rlabel metal1 83 -737 83 -737 1 p2
rlabel metal1 4 -693 4 -693 3 A2_inv
rlabel metal1 4 -781 4 -781 3 A2_inv
rlabel metal1 118 -694 118 -694 7 A2
rlabel metal1 48 -676 48 -676 5 vdd
rlabel metal1 68 -797 68 -797 1 gnd
rlabel metal1 4 -752 4 -752 3 B2_inv
rlabel metal1 118 -719 118 -719 7 B2_inv
rlabel metal1 113 -752 113 -752 1 B2
rlabel metal1 113 -782 113 -782 1 A2
rlabel metal1 142 -678 142 -678 5 vdd
rlabel metal1 142 -733 142 -733 1 gnd
rlabel metal1 169 -733 169 -733 1 gnd
rlabel metal1 169 -678 169 -678 5 vdd
rlabel metal1 139 -709 139 -709 1 A2
rlabel metal1 150 -709 150 -709 1 A2_inv
rlabel metal1 178 -711 178 -711 7 B2_inv
rlabel metal1 166 -709 166 -709 1 B2
rlabel metal1 4 -719 4 -719 3 B2
rlabel metal1 169 -528 169 -528 5 vdd
rlabel metal1 169 -583 169 -583 1 gnd
rlabel metal1 142 -583 142 -583 1 gnd
rlabel metal1 142 -528 142 -528 5 vdd
rlabel metal1 68 -647 68 -647 1 gnd
rlabel metal1 48 -526 48 -526 5 vdd
rlabel metal1 83 -587 83 -587 1 p1
rlabel metal1 4 -544 4 -544 3 A1_inv
rlabel metal1 4 -569 4 -569 3 B1
rlabel metal1 3 -602 3 -602 3 B1_inv
rlabel metal1 4 -632 4 -632 3 A1_inv
rlabel metal1 118 -544 118 -544 1 A1
rlabel metal1 118 -569 118 -569 1 B1_inv
rlabel metal1 114 -602 114 -602 1 B1
rlabel metal1 114 -632 114 -632 1 A1
rlabel metal1 139 -559 139 -559 1 A1
rlabel metal1 150 -559 150 -559 1 A1_inv
rlabel metal1 167 -559 167 -559 1 B1
rlabel metal1 177 -559 177 -559 7 B1_inv
rlabel metal1 83 -887 83 -887 1 p3
rlabel metal1 4 -843 4 -843 3 A3_inv
rlabel metal1 4 -931 4 -931 3 A3_inv
rlabel metal1 118 -844 118 -844 7 A3
rlabel metal1 48 -826 48 -826 5 vdd
rlabel metal1 68 -947 68 -947 1 gnd
rlabel metal1 4 -902 4 -902 3 B3_inv
rlabel metal1 118 -869 118 -869 7 B3_inv
rlabel metal1 113 -902 113 -902 1 B3
rlabel metal1 113 -932 113 -932 1 A3
rlabel metal1 142 -828 142 -828 5 vdd
rlabel metal1 142 -883 142 -883 1 gnd
rlabel metal1 169 -883 169 -883 1 gnd
rlabel metal1 169 -828 169 -828 5 vdd
rlabel metal1 139 -859 139 -859 1 A3
rlabel metal1 150 -859 150 -859 1 A3_inv
rlabel metal1 178 -861 178 -861 7 B3_inv
rlabel metal1 166 -859 166 -859 1 B3
rlabel metal1 4 -869 4 -869 3 B3
rlabel metal1 83 -1037 83 -1037 1 p4
rlabel metal1 4 -993 4 -993 3 A4_inv
rlabel metal1 4 -1081 4 -1081 3 A4_inv
rlabel metal1 118 -994 118 -994 7 A4
rlabel metal1 48 -976 48 -976 5 vdd
rlabel metal1 68 -1097 68 -1097 1 gnd
rlabel metal1 4 -1052 4 -1052 3 B4_inv
rlabel metal1 118 -1019 118 -1019 7 B4_inv
rlabel metal1 113 -1052 113 -1052 1 B4
rlabel metal1 113 -1082 113 -1082 1 A4
rlabel metal1 142 -978 142 -978 5 vdd
rlabel metal1 142 -1033 142 -1033 1 gnd
rlabel metal1 169 -1033 169 -1033 1 gnd
rlabel metal1 169 -978 169 -978 5 vdd
rlabel metal1 139 -1009 139 -1009 1 A4
rlabel metal1 150 -1009 150 -1009 1 A4_inv
rlabel metal1 178 -1011 178 -1011 7 B4_inv
rlabel metal1 166 -1009 166 -1009 1 B4
rlabel metal1 4 -1019 4 -1019 3 B4
rlabel metal1 282 -1018 282 -1018 1 vdd
rlabel metal1 237 -1041 237 -1041 1 A4
rlabel metal1 330 -1039 330 -1039 1 B4
rlabel metal1 290 -1037 290 -1037 1 out4_inv
rlabel metal1 308 -1055 308 -1055 1 vdd
rlabel metal1 308 -1082 308 -1082 1 gnd
rlabel metal1 316 -1065 316 -1065 1 g4
rlabel metal1 290 -1155 290 -1155 1 gnd
rlabel metal1 282 -848 282 -848 1 vdd
rlabel metal1 237 -871 237 -871 1 A3
rlabel metal1 330 -869 330 -869 1 B3
rlabel metal1 290 -867 290 -867 1 out3_inv
rlabel metal1 308 -885 308 -885 1 vdd
rlabel metal1 308 -912 308 -912 1 gnd
rlabel metal1 316 -895 316 -895 1 g3
rlabel metal1 290 -985 290 -985 1 gnd
rlabel metal1 282 -678 282 -678 1 vdd
rlabel metal1 237 -701 237 -701 1 A2
rlabel metal1 330 -699 330 -699 1 B2
rlabel metal1 290 -697 290 -697 1 out2_inv
rlabel metal1 308 -715 308 -715 1 vdd
rlabel metal1 308 -742 308 -742 1 gnd
rlabel metal1 316 -725 316 -725 1 g2
rlabel metal1 290 -815 290 -815 1 gnd
rlabel metal1 282 -508 282 -508 1 vdd
rlabel metal1 237 -531 237 -531 1 A1
rlabel metal1 330 -529 330 -529 1 B1
rlabel metal1 290 -527 290 -527 1 out1_inv
rlabel metal1 308 -545 308 -545 1 vdd
rlabel metal1 308 -572 308 -572 1 gnd
rlabel metal1 316 -555 316 -555 1 g1
rlabel metal1 290 -645 290 -645 1 gnd
rlabel metal1 526 -849 526 -849 7 c1
rlabel metal1 518 -866 518 -866 1 gnd
rlabel metal1 498 -893 498 -893 1 clk
rlabel metal1 494 -874 494 -874 1 g1
rlabel metal1 466 -825 466 -825 1 clk
rlabel metal1 500 -911 500 -911 1 gnd
rlabel metal1 508 -880 508 -880 1 n12
rlabel metal1 480 -837 480 -837 1 p1
rlabel metal1 480 -854 480 -854 1 cin
rlabel metal1 500 -850 500 -850 1 n11
rlabel metal1 509 -820 509 -820 1 vdd
rlabel metal1 626 -849 626 -849 7 c2
rlabel metal1 618 -866 618 -866 1 gnd
rlabel metal1 598 -893 598 -893 1 clk
rlabel metal1 594 -874 594 -874 1 g2
rlabel metal1 566 -825 566 -825 1 clk
rlabel metal1 600 -911 600 -911 1 gnd
rlabel metal1 608 -880 608 -880 1 n22
rlabel metal1 580 -837 580 -837 1 p2
rlabel metal1 580 -854 580 -854 1 c1
rlabel metal1 600 -850 600 -850 1 n21
rlabel metal1 609 -820 609 -820 1 vdd
rlabel metal1 726 -849 726 -849 7 c3
rlabel metal1 718 -866 718 -866 1 gnd
rlabel metal1 698 -893 698 -893 1 clk
rlabel metal1 694 -874 694 -874 1 g3
rlabel metal1 666 -825 666 -825 1 clk
rlabel metal1 700 -911 700 -911 1 gnd
rlabel metal1 708 -880 708 -880 1 n32
rlabel metal1 680 -837 680 -837 1 p3
rlabel metal1 680 -854 680 -854 1 c2
rlabel metal1 700 -850 700 -850 1 n31
rlabel metal1 709 -820 709 -820 1 vdd
rlabel metal1 826 -849 826 -849 7 cout
rlabel metal1 818 -866 818 -866 1 gnd
rlabel metal1 798 -893 798 -893 1 clk
rlabel metal1 794 -874 794 -874 1 g4
rlabel metal1 766 -825 766 -825 1 clk
rlabel metal1 800 -911 800 -911 1 gnd
rlabel metal1 808 -880 808 -880 1 n42
rlabel metal1 780 -837 780 -837 1 p4
rlabel metal1 780 -854 780 -854 1 c3
rlabel metal1 800 -850 800 -850 1 n41
rlabel metal1 809 -820 809 -820 1 vdd
<< end >>
