* SPICE3 file created from and2.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY=1.8
.option scale=1u

Vdd	vdd	gnd	'SUPPLY'
vin_x1 A 0 pulse 0 1.82 0ns 1ns 1ns 20ns 40ns
vin_x2 B 0 pulse 0 1.82 0ns 1ns 1ns 40ns 80ns

M1000 a_49_n109# A out_inv Gnd CMOSN w=10 l=2
+  ad=100 pd=60 as=50 ps=30
M1001 vdd B out_inv w_n18_n7# CMOSP w=20 l=2
+  ad=300 pd=150 as=200 ps=100
M1002 out out_inv vdd w_n18_n7# CMOSP w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1003 a_49_n109# B gnd Gnd CMOSN w=10 l=2
+  ad=0 pd=0 as=100 ps=60
M1004 vdd A out_inv w_n18_n7# CMOSP w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 out out_inv gnd Gnd CMOSN w=10 l=2
+  ad=50 pd=30 as=0 ps=0
C0 w_n18_n7# Gnd 3.84fF

.tran 0.1n 200n

.control
set hcopypscolor = 1 
set color0=white 
set color1=black 
set color2 = red        
set color3 = blue       
set color4 = green
set color5 = purple
set color6 = yellow

run
plot  v(out) v(A) v(B)
.endc